FÖRRÄDARENS LÖN

Berättelse frän sista finska kriget

Af

J. O. ÅBERG






Stockholm,
F. & G. Beijers förlag
1891.





      "Sveko vi vid Siikajokis, när det ändligt gälde se'n?"

                      RUNEBERG, Fänrikens Marknadsminne.



INNEHÅLL:


    I. Inledning. Hjertestrider.
   II. Branden.
  III. Under drabbningen.
   IV. På fädernehemmets ruiner.




I.

Inledning. Hjertestrider.


Ehuru ganska svåra strider utkämpats under det finska hären långsamt
drog sig norr ut, hade ingenting vunnits med dessa blodsutgjutelser,
annat än att den tro på ryssarnes öfverlägsenhet, som börjat göra sig
allt mera gällande bland gemenskapen, blef starkare för hvarje dag. De
exempel på feghet, som fältmarskalk Klingspor dag ut och dag in gaf
sina underlydande, kunde icke annat än uppväcka misstroende mot honom
och en dyster modstulenhet i soldaternas hjertan. De fingo ej, såsom de
önskat, och ännu önskade, på fullt allvar taga itu med den hatade
fienden; kom det någon gång till affär, och finnarne vunno någon
framgång, strax kom fältmarskalkens order om återtåg. Förbittringen och
afskyn mot Klingspor gaf sig också luft i mångahanda utgjutelser, men
hvad bekymrade det denne "kommissariatets man"; han såg endast på sin
egen fördel, och vid sitt rikligt försedda bord klagade han ändå öfver,
att han måhända skulle svälta ihjäl i Finland. Och hans soldater då,
hur lefde väl de? Illa klädda och med knapp föda måste de, genomtågande
sina fäders land såsom flyktingar, i oafbrutna strider kämpa mot en
öfvermodig, hånande fiende. Och ändå sveko de icke sina fanor. Tvärtom
strömmade nya skaror till hufvudhären, och icke nog dermed, på
landsorten erbjödo sig bönderna sjelfmant, mot det att de undfingo
gevär och ammunition, att i de vidsträckta skogarne göra fienderna allt
möjligt afbräck. Och denna glödande fosterlandskärlek, hur upptogs den
väl af "mannen med två hakor och ett öga", och af den svenska
regeringen? Det är sorgligt att påminna sig denna dystra tid, men för
att bilda sig ett rätt begrepp om detta på nederlag och härliga segrar
så rika fälttåg, måste man också se skuggsidorna.

Bönderna fingo icke de vapen, som de begärde; de blefvo tvärtom ofta
utsatta för de förnämares hån; deras ädla sjelfuppoffring betraktades
från vissa håll såsom vansinne, och om bönderna, såsom ganska ofta
inträffade, öfverraskade och nedgjorde smärre fiendtliga afdelningar,
sågs detta med visst icke blida ögon.

Siikajokiån, Sikån -- icke Sikajokiån Svinån, såsom man ibland får se
namnet stafvadt -- är omkring 400 alnar bred. Den södra stranden, på
hvilken kyrkan, prestgården, klockargården, Gerthela gästgifveri och
flere torp af betydenhet ligga, är betydligt högre än den motsatta, och
bar vid tiden för denna berättelse en ymnig skog. Ungefär 1,000 alnar
söder om kyrkan fanns en ganska djup dalgång, som man antager har
utgjort den gamla flodbädden. Bakom denna dalgång hade andra brigaden,
anförd af Georg Karl von Döbeln, intagit en fast position. På båda
sidor om vägen hade han förlagt en bataljon björneborgare, bakom midten
Österbottens södra bataljon, och bakom venstra flygeln återstoden af
björneborgarne. Vid Gerthela stodo tvenne sexpundiga kanoner. Tredje
brigaden, som utgjorde venstra flygeln af hären, hade fått sin plats på
elfvens norra strand. Andra brigaden hade redan förut blifvit afskickad
för att bemäktiga sig Carlo, en högst vigtig punkt, under närvarande
omständigheter. Adlercreutz återkallade genast denna sist nämde brigad.
Trossen, som mest varit utsatt för ryssarnes angrepp, fördes
oförtöfvadt fram på vintervägen till Sumijoki, för att alltid vara i
säkerhet.

Det var den adertonde april 1808, annandag påsk, som drabbningen vid
Siikajoki utkämpades.

Vi skrifva en af de första dagarne i april månad. Det var på
eftermiddagen, och skymningen började redan kasta sina slöjor öfver den
här och der bländhvita jorden, öfver trädens gungande snöfransar och
öfver Siikajokielfvens samt det bundna hafvets ismassa. Kölden, som de
föregående dagarne icke varit särdeles stark, hade den nämde dagen
tilltagit, hvarjemte den svaga nordanvind, som böjde trädens tunga
toppar, också bidrog till att öka kölden. Så långt blickarne kunde nå
utefter hafvet, var isfältet ödsligt, endast de der och hvar till en
ansenlig höjd upptornade islagren samt den långt i vester sig höjande
Garlön bidrogo till att något minska den enformighet, som annars skulle
vidlådt vintertaflan. Lät man blickarne deremot halka öfver den frusna
elfven, kunde det hända, att man då och då såg en enslig vandrare
skynda öfver från den ena stranden till den andra. Den tafla, som åt
detta håll upprullades för betraktarens blickar, hade icke den förras
enformighet, men öfver den låg äfven vinterns stillhet som en kylande
boja.

Vid Siikajokielfvens mynning och på dess norra strand låg ett hemman,
som vi vilja kalla Pirrtis. Det var ett af de vackraste och på samma
gång bästa som fanns i trakten, samt egdes af den högdragne bonden
Pekka Pirrtiainen. Ingen i hela trakten kunde mäta sig med honom i
egodelar; ingen kunde heller uppvisa en så väl tillredd jord som Pekka.
Detta bidrog också till att öka hans högmod, som tidt och ofta skaffade
honom stort obehag, ty de andra hemmansegarne läto icke kufva sig af
den rytande Pirrtiainen, hur väldig stämma han än hade. När denna
ovänskap först började, trodde likväl alla, att den snart skulle
upphöra och ett godt förhållande inträffa, men deruti misstogo de sig,
ty Pekka, som egentligen till sin födsel var från södra Österbotten,
och således hade dessa inbyggares olater, ville icke på några vilkor
taga första steget till försoning. Det var en styfhet utan like. Skulle
den böjas eller ej?

Det var halfmörkt i Pekka Pirrtiainens hvardagsstuga, öfver hvars här
och der bristfälliga golf han vandrade med stora steg och under det han
tidt och ofta fäktade med armarne, Pekka var mäkta upprörd, det syntes
tydligt på honom; hans små, mörka ögon glänste oftast som glimrande
eldkol, och de tunna, hopbitna läpparne tillkännagåfvo mer än tydligt,
att den kalla beräkningen, som så ofta förändrar en menniska, också
låtit honom komma på andra tankar.

"Elli tycker om honom och han om henne", mumlade Pekka och ökade
stegen. "Ja, nog är Rietu [Fredrik] bra, men han är för mycket lugn.
Ingenting förmår skrämma honom, och om faran nalkas, skrattar han henne
rakt i ansigtet. Det der retar mig, ty pojken blyges icke att skratta
äfven åt mig. _Åt mig_", fortfor han med eftertryck och knöt de
senfulla händerna. "Skratta åt mig! Nej, det skall han då inte ha gjort
ostraffadt. Rietus' far är en rysshatare af första sorten; ja, nog
hatar jag den förbannade ryssen, jag också, men", och vid dessa ord
glänste hans blickar af en besynnerlig eld, "det gör mig en ganska stor
vinst att helst vara overksam. Hvad är det för ett fördömdt påhitt, som
Rietus' far kommit upp med, att beväpna folket och i skogarne göra
fienden så mycket afbräck som möjligt! Det der lyckas aldrig, så mycket
kan jag säga, åtminstone skall jag..."

Hans monolog afbröts i detsamma, derigenom att dörren öppnades och en
ung flicka vid pass aderton år trädde in. Det var Pekka Pirrtiainens
täcka dotter, Elli, afhållen af alla och bekant för sin skönhet, äfven
långt utom Siikajoki. I det ögonblick den unga flickan trädde in, låg
ett djupt vemodigt uttryck öfver hennes drag.

"Hyvää ilta (god afton), fader", hviskade hon med en stämma, lindrigt
darrande. "Har ni hört den stora nyheten?"

"Nej, hvilken nyhet", frågade Pekka.

"Att de våra nalkas hitåt, förföljda af ryssarne?"

Hur modig Pekka än var, kunde han icke betvinga en obehaglig känsla,
som intog honom vid Ellis ord: förföljda af ryssarne. Den inre stämma,
som ropade efter mera guld, och som döfvade alla betänkligheter hos
honom, nedtystades för några ögonblick. Ellis ord kommo honom att i
dessa sekunder skåda allt det namnlösa elände, som hotade hans
fädernebygd. Men, såsom vanligt händer, de goda rörelserna voro allt
för svaga för att vinna stadigt fäste; de verldsliga bestyren togo
snart öfverhanden.

"Bah", utbrast han efter en stunds begrundande och började åter sin
vandring öfver golfvet. "Om ryssen kommer, så skall han nog uppföra sig
skonsamt; jag är säker derpå."

"Ja, lika skonsamt som öfverallt i landet, der han tågat fram", inföll
Elli, icke utan en viss bitterhet, som djupt skakade Pirrtiainen. Men
denne slog å nyo "döförat" till för det varnande i dotterns ord, och
sade i stället med allvarlig stämma:

"Du tycker om Rietu, jag vet det."

Elli spratt till. Dessa ord hade hon icke väntat sig få höra.

"Nå", sade Pekka och drog Elli fram till fönstret, på det att han
bättre skulle kunna observera uttrycket i hennes anlete, "har jag inte
rätt?"

"Jo, fader", svarade Elli sakta och lät hufvudet sjunka ned mot
bröstet. "Men", fortfor hon och upplyfte det snart, liksom insåge hon
genast, att hennes unga kärlek till Rietu icke var någonting att blygas
för, "hvarför gör ni mig denna fråga och det på ett så besynnerligt
sätt?"

"Derför, att jag icke gillar din kärlek till _honom_", svarade Pekka
med tonvigt på sista ordet.

"Hvarför då, fader?"

"Derför... derför... ah, hvad tjenar det till att upprepa det", sade
Pirrtiainen med en viss oro.

"Jo, fader, jag vill veta det", utropade Elli och omfattade lifligt
faderns arm. "Ni _måste_ säga det."

"Jaså, _måste_ jag säga det?"

"Ja."

"Nåväl då", inföll Pekka med dyster stämma, och återtog sin häftiga
gång, "Rietu och hans far stå i vägen för mina planer. Du känner dem",
fortfor han och grep Elli våldsamt i armen, "och förbannad vare du, om
du yppar ett halft ord om dem."

Elli sprang tillbaka, hennes hjerta bultade våldsamt; hon lade båda
händerna öfver bröstet liksom för att hämma de oroliga slagen.

"Nåå", utbrast Pekka dystert, "inser du inte nu, hvarför jag ogillar
din kärlek?"

"Jag kan ej upphöra att älska honom", sade Elli, icke utan
ansträngning.

"Du måste", röt Pekka till och stampade i golfvet.

"Nej, fader, jag kan icke."

"Då förskjuter jag dig och..."

"Håll", ropade Elli och sprang fram till den gamle, som dyster stod
framför henne, "vid minnet af min moder, som ni älskade så högt, besvär
jag er, att ni tager edra ord tillbaka."

"Aldrig" svarade Pekka hotande, och hans mörka ögon glödde af en hatets
eld. "Aldrig återtager jag mina ord."

En hård strid utkämpades inom Elli; det var striden om kärleken till
fadern eller till Rietu. Det blef för en stund tyst i stugan; till och
med Pekka hade slagit sig ned på en stol och öfvertänkte, med ansigtet
doldt i båda händerna, sina planer.

"Fader", sade ändtligen Elli och hennes stämma var nu fastare, "jag kan
ej svika min kärlek till Rietu, hellre..."

"Tyst, flicka", dundrade Pirrtiainen och sprang upp. "Icke ett enda ord
mer om den saken. Tyst."

Elli drog sig darrande tillbaka, ty hon visste allt för väl, att fadern
icke var att leka med, då han blef ond. Sedan hon förblifvit stum några
minuter, ämnade hon just å nyo tilltala fadern, när dörren åter rycktes
upp och en högväxt yngling inträdde.

"God afton, fader Pekka", sade Rietu, i det han skakade snön ifrån sig,
"jag har en helsning från far att tillföra eder."

Pekka mumlade för sig sjelf några ord, hvilka ej kunde förnimmas af de
andra. Härunder tog Rietu tillfället i akt att närma sig Elli och
tillhviska henne några kärlekens ord.

"Nå, hvad är det för en helsning du medför?" sade ändtligen Pekka,
sedan han en stund med kufvad harm betraktat de unga, som tycktes helt
och hållet hängifva sig åt sin kärlek. "Säg ut fort och stå inte och
prata dumheter med flickan."

En fin rodnad af förtrytelse uppsteg vid dessa Pirrtiainens skarpa ord
på Rietus kinder. Han återhöll likväl de hårda ord, som han hade på
tungan, och sade i stället:

"Ryssen nalkas. Han bränner och härjar hvar han går fram. Det är nu
fars och många andras önskan, att ni följer med, för att göra fienden
afbräck annars..."

Rietu tystnade och kastade en blick, full af smärta, på Elli, hvilkens
hjerta bultade med hårdare slag vid afhörandet af Rietus ord.

"Annars", upprepade Pekka försmädligt och satte båda händerna i
sidorna, "hvad menar du med det der ordet?"

Rietu teg en stund. Pekka upprepade sin fråga, och det nu i hotande
ton.

"Jo, annars blir ni ansedd som en förrädare." Dessa ord uttalade Rietu
lågt och med sväfvande stämma. Fruktade han måhända, att någon obehörig
lyssnare skulle finnas?

Pekka teg en stund; han kämpade synbarligen med sig sjelf en hård kamp.
Slutligen sade han med stränghet:

"Helsa du din far och alla de andra, att Pekka Pirrtiainen går sin bana
fram utan att bry sig om hvad andra tycka och göra. Du har mitt besked,
och det är att jag _icke_ följer er."

"Far, far", utbrast Elli och störtade fram till den gamle, "betänk..."

Den gamle gjorde en afvärjande rörelse med handen.

"Betänk du sjelf hvad _jag_ har sagt", afbröt han strängt.

"Ja, det har jag betänkt", svarade Elli modigt.

"Och det är?"

"Att jag följer Rietu", utbrast den unga flickan och kastade sig i
ynglingens armar. "Gud skall nog förlåta mig denna olydnad."

Uttrycket i Pekkas ansigte var hotande, och han hade den förfärliga
förbannelsen på sina läppar, men blef helt och hållet förstummad af
öfverraskning, då Rietu och Elli, utan att bekymra sig om Pekkas vrede,
störtade ut. En lång stund förgick, utan att han kunde tänka en enda
redig tanke, men slutligen återfick hans själ den spänstighet, som den
saknat under de förflutna ögonblicken.

"De ha hotat mig", utbrast han och stampade i golfvet, "men jag skall
visa dem, att Pekka Pirrtiainen alls icke fruktar deras hotelser."

Det blef nu tyst i Pekkas stuga; ingen vänlig qvinnohand ordnade såsom
förut, ty Elli hade begifvit sig till Rietus far. Hennes kärlek till
Rietu var allt för stark, att den skulle kunna rubbas. Väl tyckte hon
ibland, att hon gjorde orätt, då hon öfvergaf fadern, men hon hyste
ändock den föreställningen, att hon, på den plats hon nu var, skulle
kunna verka mera till faderns fördel, än om hon stannade qvar i hemmet,
och detta var egentligen orsaken till, att hon för ögonblicket
åsidosatte sina pligter såsom dotter. Om hon lyckades i sina ädla
bemödanden att rädda fadern, eller icke, det tillhör just denna
berättelse att lösa.




II.

Branden.


Det var påskdagsaftonen den 17 april 1808. I Siikajoki kyrkby och der
omkring rådde stor liflighet, ity att de finska bataljonerna kommit
dit. Skulle väl återtåget fortsättas längre norr ut, så frågade sig en
hvar, men han, som på denna fråga skulle svara, nemligen Klingspor, han
fanns icke vid hären. Feg som han var, hade han redan afrest mot
norden, lemnande åt Adlercreutz, som efter drabbningen vid Pyhäjoki
blifvit generaladjutant, att leda händelsernas gång. Ett hade
Klingspor, sin vana trogen, dock förständigat Adlercreutz, och det var
att genast retirera, så fort fienden envist trängde på. Det är
sorgligt, men sant: dagens lösen var detta enahanda: tillbaka! Skulle
äfven nu denna lösen utdelas?

Vi förflytta oss till en sprakande lägereld invid Siikajoki kyrkmur.
Vid elden, som flitigt underhölls, lågo tvenne björneborgska soldater
och samtalade ifrigt. Ett litet stycke ifrån dem fanns en annan bivuak,
der några officerare af olika regementen samspråkade. Och hvilket ämne
skulle väl afhandlas, om icke just kriget.

"Du, Jussi", sade den äldre soldaten och upplyfte hufvudet samt
betraktade skarpt kamraten, "har du hört, att fältmarskalken vägrat
bönderna gevär?"

"Ja, nog har jag det", svarade den, som kallades Jussi, "men jag har
också förnummit, att Siikajokis byamän sjelfve skaffat sig sådana och
för några dagar sedan tågat ut, under anförande af en bonde vid namn
Ollola. Det är käckt folk, skall jag säga."

"Ja, om det är sant."

"Jo, det är sant", inföll en underofficer, som nu trädde fram till
bivuaken; "jag hörde det för en stund sedan af dem der borta." Vid
dessa ord pekade han på officerarnes lägereld, hvarifrån ett högljudt
sorl började höras.

"Men", fortfor den gamle soldaten och reste sig upp, "det är väl inte
tänkbart, att vi få slås på allvar ännu."

"Jo, det torde allt hända", inföll underofficeren. "Både Adlercreutz
och Döbeln ha beslutat att göra skarpare motstånd här än annorstädes."

Ett tviflande leende visade sig kring den unge soldatens läppar, då han
sade:

"Deras vilja är icke gällande, såsom vi nogsamt känna till. Det är ju
Klingspor, som för befälet."

"Och som är den förste på flykten, ja", inföll underofficeren, i det
han harmfullt bet ihop tänderna.

I detsamma hördes sorlet starkare från officerarnes lägereld, och
åtskilliga utrop, sådana som "lefve Adlercreutz, lefve Döbeln",
förnummos tydligt. Inom kort var platsen mellan de båda lägereldarne
uppfyld af officerare och soldater, som uppmärksamt lyssnade till
hvad än den ene, än den andre sade. Allmänna samtalsämnet var
Siikajokiböndernas utmarsch. Jemväl spårades en tydlig oro hos alla
öfver de käcka böndernas öde, ty de hade, oaktadt fyra dagar gått till
ända, ännu icke afhörts. Hade de månne dukat under för de öfverlägsna
fienderna?

Det led allt längre och längre fram på qvällen. Skymningen öfvergick
till mörker och bivuakeldarne lyste i följd deraf klarare. Det var en
lugn och stjernklar afton, en sådan, då jorden, svept i sin hvita
oskuldsmantel, tyckes ligga försänkt i heliga böner inför all tings
upphofsman. Det var en afton egnad helt och hållet åt friden. Täflande
i hvithet med snön, låg der det åldriga templet; dess spira pekade,
såsom ännu i dag, manande upp till himmelen, och från dess torn ljöd
aftonklockans klingande toner. De manade också till frid och hvila. Men
hvad hvila kunde förunnas den på återtåg stadda hären? Kringsvärmade af
Kulneffs vaksamma kosacker, måste soldaterna i sina qvarter sofva på
geväret, beredda hvarje minut att bryta upp och genom snödrifvor och
öfver oländiga marker fortsätta det nesliga återtåget. Hvem kan då
undra på, om harmen bröt ut i ord, och det skarpa ändå; i tillmålen,
som i andra fall icke blifvit ostraffade.

Aftonklockans toner hade nyss förklingat, då en liten trupp marscherade
fram längs åns södra strand. Det syntes tydligt, att det icke var
reguliera trupper. Kanske att det var fångar.

"Der ha vi bönderna", utropade Jussi så högt, att alla kunde höra det
"Jag är säker på det."

Ett sorl af förvåning genomlopp soldathopen, ty hvar och en kunde nu
öfvertyga sig om riktigheten af den unge soldatens utsago.

Med Ollola i spetsen tågade Siikajokibönderna fram till officerarnes
bivuak. De förde med sig tio fångar, deribland en officer. Denne blef
väl mottagen och under bevakning afförd till högqvarteret.

"Ryssen är oss i hälarne", ropade Ollola.

"Det känna vi nog till", svarade en starkt byggd nyländsk jägare.

"Ja, Gud låte honom bara komma inom skotthåll", inföll en björneborgare
med stridslysten min, "nog ska vi märka honom."

"Nu till Pekka Pirrtiainen", fortfor Ollola. "Det är en förrädare och
förtjenar derför en sådans öde. Framåt, kamrater!"

"Till Pekka, till landsförrädaren Pirrtiainen!" ropade soldaterna och
bönderna om hvarandra, och öfver det döfvande larmet förnams tydligt
detta utrop:

"Tänd eld på den skurkens näste! Det förtjenar ej bättre öde."

"Ja, till Pekka!" ropade alla om hvarandra, "och låtom oss först som
sist bränna upp den skurken."

När den stora massan blir retad, är den fruktansvärd i sin vrede; den
skyr inga hinder för att nå sitt mål; den är oemotståndlig likasom
hafvets våg, som bryter öfver det redlösa fartyget.

Pekka Pirrtiainen var, såsom förut blifvit nämdt, mycket hatad af
befolkningen, icke blott i Siikajoki, utan äfven i närgränsande
socknar, och det för sin ryssvänlighets skull. Och det var naturligt,
att i denna tid, då hvarje redlig finne med gladt sinne offrade lif och
blod för fädernejordens befrielse, ett förräderi, sådant som
Pirrtiainens, icke skulle förblifva ostraffadt.

"Till Pirrtis!" ropade gamle Ollola och svängde musköten öfver sitt
hufvud.

"Till Pirrtis, till Pirrtis", skränade soldater och bönder om
hvarandra. "Död åt förrädaren!"

Det fanns en, som icke tog del i skränet, men som ovilkorligen rycktes
med strömmen. Det var Rietu. Dyster och fåordig, följde han motvilligt
bönderna; han tänkte på Elli. Ack, hur gerna skulle han icke velat
träffa henne, ty nu, då faran var öfverhängande, kände han sig manad
att bistå den skyldige, och det ehuru han var en förrädare. Rietu
tänkte icke på något annat, än att det var _Ellis_ far, som hotades af
olyckan, och att afvända denna skulle nu blifva hans förnämsta omsorg.
Men på hvad sätt skulle det gå till? Jo, endast genom att vinna tid; ty
Rietu insåg nog, att bland de församlade det allt skulle finnas någon,
som skulle underrätta Pekka om den fara, som sväfvade öfver hans
hufvud. Han sade för den skull med en stämma, som tydligt hördes af
alla:

"Låt oss vänta en stund, kanske..."

Han fick ej tala till punkt, ty en grof stämma inföll:

"Jaså, Rietu vill uppehålla oss, på det att förrädaren må kunna varnas.
Ja ja, det är inte alls underligt, när han och Elli tycka om hvarandra.
Slägten framför allt."

Rietu bleknade märkbart, och skulle just svara, då fadern utbrast:

"Perkele! Icke trodde jag mig få höra dylika ord af min son. Men är du
förrädare, pojke, du också, så känner jag dig inte, så mycket du vet
det."

Ett doft mummel genomlopp hopen vid dessa Ollolas ord, men ingen stämma
tog Rietus parti. Fanns det tilläfventyrs någon, som hyste medlidande
med den redan till döden dömde Pirrtiainen, så vågade han icke
uppträda, af fruktan för lifvet.

"Rietu håller med Pekka", hördes en stämma; "han är kanske med om
förräderiet."

"Låt oss undersöka den saken", utbrast mannen.

Då Ollola såg, att faran verkligen sväfvade öfver sonens hufvud, tog
han raskt sitt parti.

"Stilla", ropade han med dundrande stämma och höjde geväret. "Den
förste, som vågar lägga sin hand på min son, får smaka denna kula.
Rietu är ej förrädare, derpå sätter jag mitt hufvud i pant. Hvad hans
kärlek till Pirrtiainens dotter anbelangar, så är det ju en sak, som
inte rör någon af er. Framåt, kamrater! Till Pirrtis, till förrädarens
bostad!"

"Ja, ja, till Pirrtis!" ropade alla med en mun. Rietu var nu glömd;
begäret efter hämd på Pekka höll allas hjertan fängslade.

I samma ögonblick de hämdlystne bönderna och soldaterna försvunno
i skogen på norra åstranden, ilade en ung flicka, som under
öfverläggningen hållit sig dold bakom kyrkmuren och från detta
gömställe hört allt, med skyndsamma steg ned på isen. Hon tvekade några
ögonblick, om hon skulle vända om, eller icke, men slutligen tog hon
mod till sig och fortsatte sin snabba gång mot åns mynning.

"Gud låte mig ej komma för sent", flämtade hon och stannade en stund
för att hemta andan. "Gud gifve mig styrka och krafter."

Denna flicka var Elli. Målet för hennes färd gissar nog läsaren.

       *       *       *       *       *

"Far, far", ropade den unga flickan och störtade andfådd in i stugan,
"fly för Guds skull. Bönderna..."

"Hvad pratar du för dumheter", utbrast Pekka Pirrtiainen vresigt. "Lägg
dig, jag vill sofva."

"Men bönderna då", klagade Elli. "De skola mörda er, det har jag sjelf
hört."

"Hvad säger du?" sporde Pekka oroligt och reste sig till hälften upp i
sängen.

Elli omtalade i korthet hvad som förefallit vid kyrkan, och skälfvande
lyssnade Pirrtiainen derpå, ty såsom alla lömska naturer var han feg
och bar en djup förskräckelse för döden. Benen ville knappt bära honom;
hela hans kropp skälfde, som om den varit behäftad med frossan.

"Hvad säger du?" utbrast han ändtligen. "Talar du verkligen sanning?"

Elli ämnade just svara, då ett döfvande larm förnams från skogen. Far
och dotter sprungo till fönstret.

"Ja, du har rätt", mumlade Pirrtiainen med dyster stämma. "Men hvad är
att göra?" fortfor han med tydlig ångest i sina anletsdrag.

"Ni måste genast fly, fader", sade Elli brådskande.

"Och du?"

"Jag blir qvar, hvem skulle väl göra mig något illa."

"Du har rätt."

Med dessa ord grep Pekka hatten och käppen och störtade ut, följd af
Elli. Men knappt hade han tagit några steg utom dörren, då han
upptäcktes af de antågande.

"Han flyr, han flyr den skurken, den förrädaren", skreko tjogtals
röster; "hindra honom från att komma undan."

Kärleken till lifvet gaf Pekka krafter; han såg ingenting, han hörde
ingenting, utom kulorna, som hveno kring hans öron. Utåt hafvet styrde
han kosan; bland dess snöberg ville han gömma sig. Sedan jagten
fortsatts en stund, återvände bönderna med oförrättadt ärende, och
deras harm gaf sig luft i åtskilliga hårda tillmålen.

"Det är du, som hjelpt din far på flykten", sade Ollola med hotande
stämma till Elli, som i yttre dörren, till utseendet lugn, inväntade
truppen.

"Ja, det har jag", svarade Elli utan den ringaste tvekan. "Skulle ni
öfvergifvit er far, om han varit i samma belägenhet som min?"

Ollola blef svaret skyldig.

"Ja, då får flickan lida i faderns ställe", utbrast en af soldaterna.
"Hon är naturligtvis ryssvänlig, hon också."

Elli darrade. Hennes irrande blickar föllo slutligen på Rietu, hvilken,
ett rof för de djupaste sinnesrörelser, nästan vanmäktig stödde sig på
geväret. Han var nu den ende, af hvilken hon kunde hoppas hjelp.

"Nej, hon är ingen förräderska", utropade slutligen Rietu och såg sig
omkring med stadiga blickar, "och den, som vågar bära hand på henne,
han får med mig att göra. Perkele! Den som en gång till kallar henne
för ryssvänlig, han må stå sitt kast."

Med dessa ord rätade ynglingen ut sin smärta, om styrka och vighet
vittnande gestalt och intog en utmanande ställning framför Elli. Ingen
svarade på en lång stund. Ändtligen bröt gamle Ollola tystnaden med
dessa ord:

"Vi kriga ej mot värnlösa qvinnor och barn. Men Pirrtiainens stuga
skall jemnas med jorden, så mycket är säkert. Fort, gossar, tänd eld på
förrädarens näste."

Det behöfdes icke en uppmaning till. Tjogtals händer framburo
välvilligt allt, som behöfdes för att tutta på, och det dröjde icke
länge, förrän Pekka Pirrtiainens vackra gård var omgifven af ris och
qvistar.

Elli hade flytt till Rietu och snyftande hvilade hon i hans famn. Ett
svagt anskri bröt fram öfver hennes läppar, när de första eldtungorna
girigt började slicka väggarna. Snart skulle det blott återstå en
glödande askhög af det kära hemmet. Ellis mod var tillintetgjordt; hon
var å nyo den svaga qvinnan.

"Var lugn, käraste vän", tröstade Rietu och smekte den unga flickans
kinder, "det kommer väl en bättre tid."

"Men far, far", snyftade Elli. "Tänk för hvilka faror han är utsatt.
Kanske skall han frysa ihjäl, kanske blifva tagen af de otäcka
kosackerna! O, min Gud, om blott detta vore väl öfverståndet!"

Bönderna och soldaterna jublade i kapp, när eldens häftighet allt mera
tilltog. Men långt ute på hafsisen, mellan ett par väldiga snöberg,
icke långt från Carlöns strand, låg Pekka väl gömd. Han såg, att det
var hans gård, som gick upp i lågor, och hans förbittring kände inga
gränser. Men hvad ville han göra? Han måste tiga och lida och se till
på hvad sätt han skulle kunna undgå faran att falla i sina landsmäns
händer.

När Pekkas gård var något mer än till hälften nedbrunnen, dånade
larmtrumman från Pietola, och i det obestämda ljus, som snön kastade
öfver alla föremål, kunde man upptäcka mörka massor, som från det
bundna hafvet närmade sig stranden.

Det var kosackerna, som nu å nyo började den blodiga leken.




III.

Under drabbningen, i.


1.

Det var annandag påsk den 18 april 1808, som finska härens öde skulle
afgöras. Från alla håll och kanter stormade de ryska kolonnerna in på
finnarne, som enligt befallning till en början försvarade sig ganska
lamt. Adlercreutz var betänkt på att återtåga, hellre än att riskera
hären. Med dyster blick stod han på en höjd invid kyrkan, och hans ögon
öfverforo spanande allt, hvad som kom i hans väg, så väl de finska som
de ryska anstalterna. Det var vid middagstiden. Vid Pietola, der
trossen befann sig, hade Nylands jägare och dragoner mycket att göra,
och det var endast de förres ihärdiga eld, som kunde tvinga Kulneffs
kosacker att stanna. Så fortgick striden utefter hela linien, och
klockan blef ändtligen fyra på eftermiddagen. Då, sedan första och
tredje brigaden gått öfver elfven, fick Döbeln befallning att retirera.
Han gjorde det ogerna, ty den ställning, han intagit bakom den förut
nämda dalgången, gjorde, att han ansåg sig ännu längre kunna hålla
stånd. Men han måste lyda order. I den allra bästa ordning öfvergick
han för den skull isen, och stälde marschen till Karinkarda. I och med
andra brigadens återtåg fingo ryssarne större spelrum, och de ansågo
sig redan såsom herrar på platsen. En allmän stormning mot norra
stranden företogs; det såg mörkt ut för den adlercreutzska hären, ty
fienderna hade vid Grytila hemman gått öfver ån till Sadinperä, samt
hade lyckats fatta posto vid sjelfva elfvens mynning, i närheten af
Gerttula gästgifvaregård. Vi förflytta oss fram till klockan 6 på
aftonen. Den lätta skymningen hade redan inbrutit. På elfvens is och
uppför den norra stranden krälade ryssarne som i en myrstack, allt
under det finnarne med harmen i hjertat långsamt drogo norr ut. Det var
ett dystert skådespel. Mången ärrig kämpe sedan Gustaf III:s krig grät
raseriets tårar, mången tvang tåren ned igen och svor ve och
förbannelse öfver upphofsmannen till detta nesliga återtåg. Men alla
lydde, ingen vägrade att gå.

Från en liten snöhöljd kulle helt nära den plats, der von Herzen stod
med sina nyländingar, tog Adlercreutz en ytterligare öfverblick af
ställningen. Det ena smärtsamma uttrycket efter det andra vexlade i
hans manliga anlete, och mången gång frammumlade han stympade meningar,
dem ingen mer än han förstod. Han var finne till lif och själ och född
i Nyland. Det var också derför som han särdeles omhuldade krigarne från
detta landskap. Framför honom låg det öfvergifna Finland, prisgifvet åt
den härjande fienden; bakom honom den höga, kalla norden med sin is och
sin snö; omkring honom hans pröfvade soldater, färdiga att lida,
färdiga att kämpa till sista man. Hvad skulle han icke tänka i dessa
ögonblick; hur smärtsamt skulle icke hjertat krympa tillsammans vid
tanken på det kommande! Adlercreutz for med afviga handen öfver den
svettiga pannan, och en djup suck banade sig väg ur hans bröst. Hans
blickar föllo på nyländingarne, och de ljusnade en smula. Hans
forskande öga mötte von Herzens. Var det måhända denna blick som med
ens förändrade stridens gång?

Ryssarne trängde på, och minut efter minut blef finnarnes trångmål
större. Då sprängde Adlercreutz på sin eldiga springare fram till von
Herzen. Hans öga brann af feberns glöd och hans stämma darrade
lindrigt, då han utropade: "Tillbaka!"

Von Herzen rörde sig ej; hans soldater stodo likaledes orörliga som
bildstoder.

Adlercreutz studsade; detta hade han icke väntat sig. En skär rodnad
sprang upp på hans kinder, och han var nära att förifra sig.

"Tillbaka", ropade han med stränghet, och det blanka svärdet blänkte i
hans hand.

Von Herzen kastade en pröfvande blick öfver sina tätt sammanslutna led.
Det brann äfven i hans ögon en flammande eld; hans hjerta bultade
våldsamt och hans senfulla hand omfattade konvulsiviskt svärdfästet.

"Tillbaka, tillbaka", dundrade Adlercreutz med hotfull stämma.

Då sprang von Herzen fram i têten af sin kolonn; hans kinder brunno som
af feberns eld, hans blickar tycktes genomborra hvarje soldat, och hans
väldiga stämma lät som åskan, då han, höjande svärdet öfver sitt
hufvud, ropade:

"Framåt! fäll bajonett!"

Nu blef det lif i den förut till utseendet stendöda kolonnen; ett
enstämmigt utrop af glädje förnams; bajonetterna fäldes så fort som de
kanske aldrig förut blifvit fälda; den jemna marschen ökades med hvarje
sekund, och många minuter hade icke gått till ända, då kolonnen med
stormsteg rusade nedför stranden, öfverändakastande allt i sin väg.

Adlercreutz visste knappt till sig, han rycktes med i strömmen; hans
entusiasm lågade å nyo upp; hans springare var som af eld, och sjelf i
spetsen för de modiga nyländingarne, högg han in på de ryska
kolonnerna, som vacklade, dels krossades, dels förströddes som agnar
för vinden.

"Löjtnant", ropade han till sin adjutant under sjelfva stormningen af
södra stranden, "spräng å stad; kalla de andra brigaderna tillbaka. Vår
är segern!"

Herzens bataljon hade, lik en lavin, med oemotståndlig makt sprängt
ryska centern. Blod och död betecknade dess väg. Nu blef det annat af.
Från alla håll återkommo de finska afdelningarna. Trögt hade de tågat
tillbaka; nästan i språngmarsch vände de åter. Ack, deras heligaste
önskan, att få på fullt allvar mäta sig med den hatade fienden, den
skulle nu uppfyllas, de skulle få visa, att de hade mod i bröstet och
kraft i armen. Hvilket ändlöst jubel, när de vikande massorna kastade
sig öfver fienden; hvilken ryslig förvirring; hur stolt och segerglad
ljöd icke björneborgsmarschen öfver stridsbullret; det var ett helt
folk, smädadt, tillbakasatt, jagadt nära nog ur dess landamären, som nu
i ett ögonblick fick vakna upp till en annan verklighet, i hvilken
segerns krona vinkade så skön; det var en berusning, som var omätlig;
om mångdubbel styrka stått emot dem, skulle finnarne ändå vunnit seger.

Då centern så oförmodadt genombröts, måste de båda ryska flyglarne, som
just höllo på att förfölja den finska hären, retirera, för att icke i
sin ordning blifva öfverflyglade. Det dröjde icke länge, förrän striden
å nyo utspann sig längs hela norra stranden, upp på hvilken ryssarne
blifvit jagade, snart sagdt i en handvändning.

       *       *       *       *       *

Dyster och ett rof för de gräsligaste lidanden vandrade Pekka
Pirrtiainen mellan de kylande snöbergen. Fram till Siikajoki tordes han
icke. Förrädarens samvetsförebråelser hopade sig öfver honom och tyngde
hans sinne; hvart han såg, tyckte han sig upptäcka armar, som ville
gripa honom, krossa honom. Under det Pirrtiainen fridlös irrade
omkring, hade Rietu slutit sig till en ströfkår, som blifvit utsänd för
att undersöka isen. Den unge mannen brann af begär lika mycket att
utmärka sig, som att få reda på Pekkas spår. Och detta för Ellis skull.

Det var stark skymning, då den trupp, till hvilken Rietu hörde, tågade
ut i riktning mot Carlön. Truppen var sammansatt af nyländingar och
björneborgare; hvar och en täflade att göra sitt bästa; här och der
skingrades en trupp ryssar, här och der tillfångatogs en annan. Elden
från handgevärssalvorna upplyste de kala snödrifvorna och spred ett
magiskt, fastän minutligt sken öfver det vidsträckta, ödsliga fältet.
Ljudet från kanonerna och musköterna vid Siikajoki hördes än doft, än
klart och tydligt.

Plötsligt spratt Rietu, som gick i främsta ledet, till. Hvad kunde
orsaken vara? Jo, mellan ett par höga snödrifvor hade hans skarpa öga
upptäckt en manlig varelse, som bemödade sig om att så fort som möjligt
fly undan. Väl kunde han icke upptäcka den flyendes anletsdrag, men en
inre stämma sade honom, att det var Pekka, och han uppbjöd allt, hvad i
hans förmåga stod, att följa hans spår.

Äfven Pekka hade igenkänt finnarne. Hade det varit ryssar, skulle han
icke ett enda ögonblick tvekat hvad han borde göra: bättre att
öfverlemna sig åt fienden, än åt de förbittrade socknemännen, ty i
senare fallet visste han nog, att hans död var gifven.

Den starka kölden hade ännu icke förmått att stelna hans lemmar; det
var den inre starka spänningen, som höll hans lifliga själ i en orolig
verksamhet, som gjorde, att han icke så snart erfor köldens inverkan.

Från drifva till drifva ilade han undan allt hvad han kunde, men
finnarne voro honom städse i hälarne. Seg som en äkta österbottning,
höll han ut i det längsta, men det var dock tydligt, att, huru härdade
hans senor än voro, han ändtligen skulle duka under för tröttheten. Med
förfäran tänkte Pekka på det ögonblick, då han måste gifva sig fången.
Han gaf till ett ilsket vrålande och de senfulla händerna knöto sig
konvulsiviskt om skaftet på en bredbladig, skarpslipad knif, hvilken
han i brådskan icke glömt att taga med sig. Skulle han ännu göra ett
försök att fly undan, eller skulle han försvara sig. Han var en stund
riktigt obeslutsam om hvad han skulle företaga. Men då han ändtligen
hade beslutat sig för något och skulle begifva sig af mellan ett par
drifvor, hejdades han plötsligt af en person, som stängde hans väg.

"Ha, fader Pekka", sade Rietu och uträckte sin hand, "ändtligen har jag
funnit er. Nu skall ni icke irra omkring här längre. Döden skulle hinna
er förr eller senare."

"Låt mig gå, Rietu", bad Pirrtiainen med ångestfull stämma.

"Nej, fader Pekka, ni måste stanna."

"Du får alla mina egodelar, ja, du får Elli på köpet."

"Ni får ej gå", svarade Rietu å nyo med allvarsam stämma.

"Nej", utbrast Pekka och hans ögon glödde af en hemsk eld, "hellre
stupar jag här."

Med dessa ord svingade Pekka den skarpslipade knifven öfver sitt
hufvud. Han syntes beslutsam.

Rietu sprang fram, just som Pekka Pirrtiainen slungade en björneborgare
till marken. Utan att länge betänka sig rusade han på den gamle bonden
och slog sina armar kring hans kropp. Förgäfves ansträngde sig den
gamle af alla krafter för att slippa lös; han satt som i ett skrufstäd.

"Släpp mig", ropade han med vansinne, "jag måste blifva fri."

"Nej", svarade Rietu allvarligt; "ni måste följa mig. Jag ansvarar för
er säkerhet."

Pekka såg en stund tvinande på Rietu; dennes förklaring, att han skulle
ansvara för honom (Pekka) susade så besynnerligt i hans öron. Skulle
han, som var stämplad såsom förrädare, kunna hoppas på tillgift! Det
såg åtminstone i det närvarande mörkt ut.

"Ni måste foga er i ert öde", sade Rietu, när de öfriga finnarne
omringade dem.

"Hvar är Elli?"

"Ah, hon är i godt förvar; på henne går det rakt ingen nöd."

Detta tycktes någorlunda återgifva Pekka det lugn, han så väl behöfde.
Med en djup suck fogade han sig i det närvarande oundvikliga.

Sedan recognosceringen var fullbordad, återvände den lilla truppen till
Siikajoki och hann fram under det striden ännu pågick som bäst.


2.

Ellis sinnesstämning kan hvar och en med lätthet fatta. Visserligen
omhuldades hon på det omsorgsfullaste af Rietus mor, men det var ändå
icke detsamma: hon saknade allt för mycket den älskade, hvarjemte oron
öfver faderns öde ständigt höll hennes själ i spänning. Men Elli var en
modig och förståndig flicka, som, efter ett kort resonnemang med sig
sjelf, kom till den förnuftiga slutsatsen, att det alls icke tjenade
till någonting att sörja i otid, utan fastmera handla så långt
omständigheterna det medgåfvo. Det första, hon då bråkade sin hjerna
med, var att utfundera ett sätt att rädda fadern, i fall han, såsom hon
förmodade, skulle blifva tillfångatagen. Väl tänkte hon i vissa
ögonblick på att uppdaga allt för Adlercreutz, och hon var nära deran,
då hon en gång mötte honom, men inom hennes bröst fanns det ändock
_något_, som höll henne tillbaka. Detta något, som obevekligt stälde
sig emellan henne och lyckan, det var den omständigheten, att fadern
var en fosterlandsförrädare. Så modig Elli än var, skälfde likväl
hennes kropp af fruktan, då hon tänkte derpå.

Nu, då striden rasade som värst, skulle hon då gitta i overksamhet och
åse huru hennes bröder lemlästades? Nej, dertill var hon för mycket
qvinna, för mycket finska. Hon begaf sig ut. Visserligen studsade hon
för några ögonblick tillbaka, när kulorna började hvina omkring öronen,
men hon tog snart mod till sig, och det varade icke länge, förrän hon
var ifrigt sysselsatt med att förbinda de sårade och skaffa nödig
hjelp, så väl åt vän som fiende. Den unga flickans modiga uppträdande
aftvådde icke allenast den mörka fläck, som faderns nedriga handling
satt på henne -- hennes älskliga och milda väsende, detsamma äfven i
faran, uppväckte allas beundran, både officerares och manskaps.

"Bra gjordt, flicka", ropade en högre officer, då Elli med anlitande af
alla sina krafter drog en sårad krigare till ett af dikena och der
började bispringa honom med all den hjelp, hon för närvarande kunde
åstadkomma.

"Bra, bra", ropade flere röster bredvid den unga flickan, som,
uppmuntrad af bifallen, arbetade med den mest spända ifver. "Om alla
vore så modiga som du, skulle inte så många dö undan."

När ingenting mer var att göra på norra stranden, sprang Elli fram till
den södra, der Herzens bataljon som bäst höll på att storma. Här tyckte
den unga flickan visserligen, att det kändes ännu värre än på den andra
stranden, men begäret att utmärka sig hade så intagit henne, att det
tycktes henne vara en af de största njutningar att nu å nyo få kasta
sig in i stridsbullret. Utan betänkande följde hon de eftersta leden af
Nylands infanteri, men plötsligt stannade hon och hela hennes kropp
skälfde. Hvad såg hon månne, som så upprörde henne?

Icke så särdeles många alnar ifrån henne hade Adlercreutz för några
minuter hållit stilla och betraktade från sin farliga ståndpunkt den
sig allt mera utspinnande striden. Omkring sig hade han nu endast några
få soldater och en adjutant. Elli kunde icke taga sina vackra blickar
ifrån befälhafvaren, som satt der på sin eldiga springare, till
utseendet fullkomligt lugn, men till sitt inre ej olik en glödande
vulkan. Hvad beundrade hon hos honom? Var det väl hans uttrycksfulla
ansigte, hans väl växta kropp? Nej, hon beundrade det mod, som han
ådagalade, när han tvärt emot order bjöd fienden spetsen.

Plötsligt höjdes ett gemensamt rop af de omkring befälhafvaren varande
soldaterna, och det var äfven hög tid för Adlercreutz att sätta sig i
försvarstillstånd, ty i sporrstreck närmade sig nu en liten kosacktrupp
med dragna sablar; den styrde kosan mot Adlercreutz. Snart kom striden
äfven här i gång, och den blef ytterst hårdnackad.

Adlercreutz och hans män kämpade med verkligt dödsförakt, ty i förstone
såg det verkligen mörkt ut för dem att komma undan, alldenstund
fiendernas antal efter hand ökades, hvaremot finnarnes minskades. Kalla
till sig förstärkning ville han icke, ty då skulle måhända slagets öde
berott derpå.

"Låtom oss genombryta fiendernas led", ropade han i stället och
sporrade hästen mot den till utseendet svagaste punkten. Men då han här
mötte ett det ihärdigaste motstånd, såg han sig tvungen att afstå från
hvarje försök.

"Detta ser ut att blifva vår sista strid här på jorden", sade han till
sin adjutant, löjtnant Lange. Men denne svarade frimodigt:

"Åhnej, herr general, ännu skola vi lägga i dagen vår kärlek till vår
födelsebygd."

"Det skola vi, om vi också skola stupa derför", sade en annan af
officerarne och uppträdde vid dessa ord en svartmuskig kosack på sin
värja som en stek på ett spett.

Från Herzens bataljon hördes dånande hurrarop; den hade fullständigt
sprängt ryssarnes center; icke långt derifrån slogos björneborgarne med
ursinnig tapperhet, och lik en mörk, med en oundviklig död hotande
lavin skred den tavastländska bataljonen med Gripenberg i spetsen södra
stranden utför. Öfver Siikajokiån och de närmaste skogspartierna
simmade den qväfvande krutröken och gjorde tillsammans med skymningen
det till slut ganska svårt att igenkänna hvarandra.

Utan att Elli visste af det, hade hon, tillika med ett par andra lika
behjertade qvinnor, blifvit indragen i den hvirfvel, som omslöt den
stridande Adlercreutz. Hennes hjerta bultade våldsamt, och hennes späda
fingrar omfattade konvulsiviskt kolfven på en skarpladdad ryttarpistol,
tillhörande en fallen kosack, att döma af inskriften, hvilken den unga
flickan icke förmådde tyda. Skärande kontrast! Med ena handen höll hon
pistolen, i hvarje minut färdig att utsända den dödande kulan; med den
andra handen aftorkade hon varsamt det ymniga blod, som flöt ur en
soldats genomstungna bröst. Hon såg en kosack rikta lansen mot
Adlercreutz's bröst, musklerna i hennes arm spändes hårdare; sakta
reste hon sig från den knäböjande ställning hon intagit; i det döfvande
vimlet, der hästar, menniskor och döda föremål syntes som ett enda
kaos, en fantastisk sammangyttring, såg Elli, den modiga bondflickan
från Siikajoki, endast den fara, som sväfvade öfver generalens hufvud.
Hon bekymrade sig icke om de stridandes buller, om de sårades och
döendes qväfda utrop. Modigt och utan att darra utsträckte hon högra
armen, under det hon stödde den venstra mot en döende hästs länd. I
detta ögonblick rörde sig ingen muskel i hennes täcka anlete.

Kosacken kom närmare; de omkring Adlercreutz varande slöto sig tätare
tillsammans, hvar och en beredd att offra ända till sista blodsdroppen
för befälhafvarens räddning. Då, just i det kritiska ögonblicket,
smälde ett skott från sidan; kosacken släppte lansen; fötterna, med
hvilka han, enligt detta steppfolks vana, styrt springaren, släppte
sitt fäste; armarne beskrefvo några våglinier i tomma luften, liksom
ville de åter gripa efter vapnet; ett svagt stönande hördes från
steppsonens läppar, derpå föll han tungt till marken. De öfriga
kosackerna studsade, och detta gaf finnarne tid att å nyo samla sig och
anfalla med fördubblade krafter. Deras angrepp blef nu oemotståndligt,
och de skyndade sig undan så mycket fortare, som Kulneffs ryttarskaror
ute på hafvet nu måste jaga tillbaka, medan de finska brigaderna
erhållit befallning att vända om. Det var ett egendomligt och tillika
fängslande skådespel, att i den lätta skymningen se de ryska
kavalleriskarorna spränga öfver isen och det bländhvita snötäcket. Hade
ej kanondundret, handgevärssalvorna och de stridandes döfvande larm
tryckt sin verklighetsstämpel på taflan, skulle man trott, att allt
endast var ett fantasispel.

När de ryska massorna allmänt veko tillbaka och segern ansågs med
säkerhet vunnen, kom general Adlercreutz fram till Elli, som ännu
outtröttligt höll på att egna sårade vänner och fiender sina ömma
omsorger. Generalens ögon uttryckte en allt för tydlig beundran, och
han sade, i det han vänligt klappade den djupt rodnande Elli, som vid
hans ankomst stigit upp:

"Du har räddat mitt lif, flicka. Hvad heter du, och hvarifrån är du?"

Elli sade sitt namn och boningsort.

"Således husvill i detta krigets elände och i denna köld", mumlade
Adlercreutz halfhögt för sig sjelf. "Stackars flicka!"

Elli hade, utan att hon behöfde anstränga sina hörselorganer, förnummit
generalens ord.

"Ah, med mig är det alls ingen fara", utbrast hon och såg sig omkring.
"Jag har nog i kyrkbyn vänner, som inte skola neka mig tak öfver
hufvudet." Och med dessa ord lät hon sina blickar öfverfara några
qvinnor, hvilka, liksom hon, voro ifrigt sysselsatta med de sårade.
Dessa qvinnor förstodo mer än tydligt Ellis blickar, och i deras tysta
nickningar kunde man läsa detta: Vi äro beredda att uppoffra allt för
dig.

Detta tysta, men vältaliga språk förstod synbarligen äfven Adlercreutz,
ty han sade till Elli, i det han åter steg till häst:

"Jag ser, att du är i goda händer. Vill du utbedja dig någonting af
mig, så uppsök mig och jag skall göra allt hvad jag kan för dig."

Med dessa ord gaf talaren hästen sporrarne och försvann i stridsvimlet.

"Ja, det torde kanske snart behöfvas, att jag anlitar hans hjelp",
tänkte Elli för sig sjelf. "Det beror på, huru det går med far. Ah, nu
skall det allt gå bra", utbrast hon med inre hänförelse; "han såg ju så
mildt på mig, då han sade, att jag skulle uppsöka honom. Ja, far skall
blifva räddad, och det genom mitt lyckliga skott."

Hur lätt hoppas icke barnet och ynglingen, att allt skall utfalla efter
deras önskan; och om detta lifliga hopp ej funnes, hvad skulle då
verlden vara? Ett hemvist för själar, utan detta aningens och hoppets
sälla rosenskimmer, som mången gång förmår att nedbryta det oblida
ödets skrankor.

Då Adlercreutz lemnade Elli, hördes de första svaga tonerna från
björneborgsmarschen i södra strandens skog. Dessa toner kommo närmare;
de brusade mäktiga som åskor, och de hänförde äfven de redan i striden
stående. Den trötte kände ny kraft tillströmma armen, den sårade
ansträngde sig för att resa sig upp en smula, och kring de läppar, som
redan började skälfva af dödens kalla kyss, spred sig ett sekundlikt
leende. Ack, hvad skulle icke dessa käcka krigare känna i dessa
stunder, på denna deras första högtidsdag! Dödens smärta blef ljuf, ty
de visste att segern var deras.

Adlercreutz sprängde emot Döbeln; deras blickar möttes, deras händer
slöto sig i hvarandra. Hvad skulle icke _de_ känna i denna stund! När
de sist sågo hvarandra, fördystrade tanken på det hopplösa återtåget
deras blickar; nu deremot, nu vinkade något helt annat: den första
härliga segern.

Björneborgarne störtade som rasande lejon utför södra stranden, öfver
isen och uppför den norra stranden. Hvad de förut gående skarorna icke
kunnat drifva undan, det mejades nu som säd till marken, så vida det
icke flydde. Förgäfves förde Rajewsky och Kulneff sina skaror i elden;
de kastades öfver ända snart sagdt i en handvändning; allt måste fly,
och allt flydde.

Sådan var aftonen af annandag påsk 1808. Den utmattade här, som
tillförne måst draga sig tillbaka, hade nu rest sig upp och aftvått
skammen med en lysande seger -- en seger, som återgaf den förtröstan
till nya framgångar och gjorde fiendens tro, att han var oemotståndlig,
om intet.

Och han, som egentligen var satt till öfverbefälhafvare för den
svensk-finska hären, var han, _fältmarskalken_ Klingspor, månne
närvarande vid drabbningen och ledde dess gång? Nej; redan långt förr
än de första skotten föllo, hade han i en beqväm släde skyndat norr ut.
Han var för mycket rädd om sin värda person, att han skulle gifva den
till pris i en kamp på lif och död.

Och åt en sådan fältherre, om hvilken den genomhederlige gamle Lode i
Franzila hade det mustiga yttrandet, att

    "det är skam att tappre männer
    täckas tala om en sådan",

hade Sveriges konung och råd anförtrott försvaret af brödralandet öster
om Bottnen. Man kan icke, vid kännedomen härom, annat än erfara djupt
vemodiga känslor af en harm, som utgången af fälttåget visade vara
fullt berättigade.

En lycka var, att hären egde så dugliga och beslutsamma
underbefälhafvare som Adlercreutz, Döbeln och Sandels, annars hade
armén väl icke fått stanna förr än vid nordpolen.




IV.

På fädernehemmets ruiner.


Det var ett par timmar efter det striden ändat; finnarnes segersånger
hördes då och då genomtona luften, alla försakelser voro nu förgätna,
framför Finlands käcka söner låg nu fosterlandet å nyo öppet; den
första segern var vunnen, och långt i söder ströfvade de ryska
bataljonerna för att hinna undan i tid. Den finne, som kunde öfverlemna
sig åt sömnen, han gjorde det nu med all trygghet; den som icke kunde
det, och många voro de, ströfvade omkring på det af tusendes blod
fuktade bataljfältet, kanske för att söka en kamrat, måhända också för
att i ensamheten påminna sig de näst föregående timmarnes faror och
värma sin själ vid hågkomsten af de utkämpade bragderna.

Bland dem, som med skyndsamma steg ilade vester ut, finna vi Elli
alldeles ensam. När striden afstannat, blef det henne för trångt inom
Ollolas stuga; hon måste hemta frisk luft; hon måste, kosta hvad som
helst, ännu en gång återse det brända fädernehemmet, der hon lidit så
mycket, njutit så mycket. Det dröjde icke länge, förrän hon var framme
vid Pirrtis ruiner, från hvilka ännu en svag hvitgrå rök uppsteg mot
vårhimmelen. En dyster bäfvan genomfor den unga flickans kropp, när hon
satte foten på en af de kolade bjelkarne; hon ville ännu icke riktigt
tro, att det hon såg var den nakna verkligheten; hon gnuggade sig
häftigt i ögonen. Kanske att allt var en sorglig dröm, påskickad henne
till pröfning! Ack, nej; verkligheten var allt för sann; den kolade
bjelken knastrade under Ellis fötter, och hur mycket hon än gnuggade
ögonen, såg hon ändock, att röken alls icke var någon bedräglig
synvilla.

"O, min Gud, min Gud", suckade hon och knäppte händerna bedjande
tillsammans öfver bröstet, "det är då en ryslig sanning, att jag ej
mera har något fädernehem! Och du, min stackars far, hvar är du nu?
Kanske irrar du omkring ute på det vida hafvet och vågar dig ej fram
till bebyggda ställen!"

Vid dessa ord sprang hon upp från sin ödmjukt knäböjande ställning;
hennes ögon voro fuktiga, hennes barm häfde sig med våldsamma slag. Hon
tänkte öfver, antingen hon skulle vända om till Ollolas gård eller
begifva sig ut på isen, för att uppsöka fadern. Men nu kunde hon icke
besluta sig så fort som hon annars brukade; det var inom henne
någonting, som alltid höll tillbaka, då hon trodde sig ha fattat
beslutet.

De tunga skyarne delade sig efter hand, och Elli hade icke lång stund
varit på ruinerna, då hon omgöts af månens klara strålar. På strid
följer frid. Lugnet i naturen återgaf den unga flickan också i viss mån
lugnet i själen. Hon gick med varsamma steg öfverallt i det nedbrända
hemmet; hon undersökte allt hvad som kunde vidröras utan att falla till
stoft, och hon hade just slutat sin vandring, samt öfvertänkte nu på
nytt, hvart hon skulle styra sina steg, då ett buller, som med hvarje
minut tilltog, tog hennes uppmärksamhet i anspråk.

"Kan det vara ryssar", tänkte hon och darrade. "Nej, de äro ju slagna.
Då är det finnar. Tänk om..."

Hon fick ej tala till punkt, ty en liten trupp, som med långsamma steg
bröt fram ur strandskogen och satte marschen på Pirrtis, hejdade henne.
Truppen närmade sig; Elli gaf till ett anskri af smärta, ty i första
ledet igenkände hon fadern med bakbundna armar. Nästan medvetslös
vacklade hon fram, men hade icke uttagit många steg, förrän hon sjönk i
Rietus armar. Hennes kinder hade snöns färg, hennes läppar voro som
förseglade; hon kunde i detta ögonblick icke ens tänka redigt; en kort
vanmakt öfverföll henne. -- -- --

       *       *       *       *       *

"Mine herrar", sade Adlercrentz ungefär vid samma tid som mötet på
hemmets ruiner egde rum, till sina underbefälhafvare, och gick med
häftiga steg fram och tillbaka i det rum han tagit i besittning, "vår
ställning är nu så mycket bättre, att vi kunna gå anfallsvis till väga.
Och vi skola ej lemna tillfället obegagnadt; det återkommer måhända
aldrig mera. Nästa dust blifver..."

Ett buller utanför dörren gjorde, att han afbröt sitt tal. Han syntes
en smula missnöjd.

"Hvem är det", sporde han posten, som nu inträdde.

"En ung flicka, herr general, en ung..."

"Har synbarligen förvridit hjernan på dig", afbröt Adlercreutz tvärt
den stammande soldaten, och det med en viss skämtsam ton. "För in
flickan!"

När dörren öppnades för andra gången, var det Elli som trädde in. Snöns
blekhet hvilade ännu öfver kinderna, blickarne stirrade utan återvändo
åt alla sidor.

"Hvad vill du, flicka?" sporde Adlercreutz medlidsamt och tog Ellis
händer mellan sina. "Du är så upprörd."

Det vänliga tilltalet hade ett afgörande inflytande på Elli. Hon
lösryckte händerna, for med dem öfver pannan och tycktes en stund
öfvertänka hvad hon skulle säga.

"Tala fritt", sade generalen med en stämma så mild, att Elli spratt upp
ur sina drömmar och med ett lätt, ett gladt utrop kastade sig till hans
fötter, under det hon utropade:

"Ni förlåter ju ett brott! O, ja, jag ser det på er, general! Min far
är brottslig; han hålles för en förrädare derför, att han icke ville
följa bönderna på deras ströftåg. Vårt hem är uppbrändt, och nu vilja
Siikajoki byamän taga lifvet af min far, som lyckats fly undan, men
blifvit fångad nära Carlön. General", fortfor den vackra flickan och
sträckte bedjande sina händer mot Adlercreutz, som, sjelf ett rof för
de mest olikartade sinnesrörelser, knappast visste hvad han skulle
tänka, "ni lofvade, att jag skulle få utbedja mig någonting af eder
derför att jag räddat _ert_ lif; nu beder jag om _min fars_ lif. O,
skynda er, annars kommer ni för sent! Skynda er!"

Adlercreutz lät sina blickar en stund hvila på krigskamraterna. I
somligas ögon läste han det obevekliga svaret: "låt förrädaren undfå
sin förtjenta lön", i andras deremot, och, vi tillstå det, i de
flestas: "låt denna gång nåd gå för rätt."

"Din far skall blifva fri", sade ändtligen generalen och tecknade några
ord på en papperslapp, gaf den åt en af sina adjutanter och befalde
honom att följa Elli.

Den unga flickans glädje var outsäglig. Hon hade ju räddat sin far, och
hon var säker på, att han efter den dagen skulle börja ett annat lif.
Adjutanten kunde endast med ansträngning följa henne; lik en jagad hind
ilade hon öfver snöfälten mot fädernehemmets ruiner.

Knappt hade hon försvunnit från generalens bostad, när Adlercreutz
vände sig till de församlade, i det han sade:

"Mine herrar, det lyster mig högligen att se utgången på denna sak. Det
torde hända, att bönderna här tillämpa den grymma lynchlagen. Viljen I
följa mig?"

Alla voro genast färdiga, helst som natten var obeskrifligt härlig, och
snart voro de på väg till Pirrtis.

       *       *       *       *       *

Läsaren fattar nogsamt orsaken till Ellis plötsliga uppträdande hos
Adlercreutz. Bönderna svuro enhälligt, och med dem soldaterna, att
landsförrädaren, hända hvad som hända ville, skulle hänga i det
närmaste trädet invid sin egen sköflade gård. Förgäfves bad Elli om
tillgift för fadern, förgäfves lofvade denne att bättra sig, och lika
förgäfves tiggde Rietu om Pekka Pirrtiainens lif.

"Han måste dö", skränade bönderna och soldaterna om hvarandra.

En djup suck höjde Pekkas bröst. Han ville tala, men orden fastnade i
halsen. Det var förfärliga stunder för den fordom så högmodige bonden.
Döden gapade mot honom; endast ett underverk kunde rädda honom, det
insåg han mer än väl. Men Pekka Pirrtiainen trodde icke på några
underverk, derför underkastade han sig, åtminstone till utseendet, det
öde, som väntade honom. I hans bröst stormade dock de våldsammaste
lidelser; han måste anlita hela sin själsstyrka för att visa sig
någorlunda lugn, ty han visste, att endast detta kunde stämma hans
fiender till hans förmån.

När Elli märkte det fåfänga i att slösa med böner, delgaf hon Rietu
sitt fasta beslut att skynda till Adlercreutz, samt omtalade orsaken
till de gynsamma förhoppningar hon hyste.

"Gå du, käraste vän", hviskade Rietu; "jag skall emellertid försöka att
uppehålla bönderna och soldaterna i det längsta."

En tacksam, kärleksfull blick, och Elli var försvunnen.

Det blef en stund tyst vid ruinerna, öfver hvilka månen göt sitt bleka,
dallrande sken. Stunden var icke utan sin stora högtidlighet. Man såg
här ett folk i beredskap att hämnas på den, som med stolt förakt
trampat fosterlandskärleken under fötterna. Det var grymt, men
rättvist. Ren och stark lågade denna kärlek i österbottningarnes bröst;
de kunde icke ens tåla _höra_ namnet landsförrädare, och när dertill
kom, att den brottslige var från samma provins, ja, till och med var
bosatt i samma socken, blef hatet mot honom ännu mera uppjagadt.

En half timme hade gått till ända, och ännu hade ingen arm höjt sig för
att verkställa den redan afkunnade domen. Ville Pekkas domare grymt
leka med honom, såsom katten med råttan? Det är svårt att säga, men
skenet hade det likväl för sig.

Plötsligt utbrast en af soldaterna så högt, att det hördes öfver hela
samlingen:

"Nu tycker jag det är tid att gifva förrädaren Pekka Pirrtiainen den
lön han förtjenat."

Bönderna och soldaterna rusade upp. Äfven Rietu, som redan från början
tagit plats bredvid den lifdömde, reste sig upp och intog en hotande
ställning framför Pirrtiainen. Ynglingens ansigte var dödsblekt, och
beslutsamheten stod tydligt att läsa så väl i hans ögon som i alla hans
drag.

"Gå bort ifrån honom", röt en jättelik bonde och armbågade sig fram.
"Vi måste taga hans lif."

"Nej", utbrast Rietu med styrka, "jag lemnar icke Pekka, förrän ni
lofvat mig att ej göra honom något ondt."

"Men, betänk då, Rietu", frampustade Pirrtiainen, under det
ångestsvetten rann utför hans panna, "du utsätter ju äfven dig för
misstankar, och hvem vet hvilken hämd som..."

"Tyst, fader Pekka", afbröt den käcke Rietu beslutsamt; "endast öfver
mitt lik skola de komma er på lifvet."

"Vettvilling", skrek en medelålders bonde och sprang fram till Rietu
samt grep honom i armen, "ser du då inte, att äfven du går din
undergång till mötes, om du längre envisas att försvara förrädaren!"

"Tillgif honom då hans brott, såsom en rättvis och barmhertig Gud också
skall tillgifva honom det", bad Rietu bevekande.

"Nej", ropade alla med en mun. "Häng förrädaren!"

Pekka Pirrtiainens kropp skakades som af en frossa. Han såg nu, att
något medlidande icke stod att erhålla.

"Nåd, nåd!" stönade Pekka med skälfvande stämma.

"Nej", skreko alla om hvarandra, "upp i trädet med honom!"

"Tillbaka", dundrade Rietu och kastade en bonde till marken, samt gaf
en annan ett så häftigt knytnäfslag för bröstet, att han ryggade
tillbaka. "Endast öfver mitt lik skola ni komma till Pekka."

Det var ett egendomligt skådespel, som nu uppfördes vid Pirrtis ruiner.
Hufvudfiguren, Pekka Pirrtiainen, med dödsångsten tecknad i sina mörka
drag och skälfvande son om han legat i frossa; Rietu stående framför
honom och med de senfulla händerna höjda till slag, samt den fasta
beslutsamhet, som icke låter rubba sig af någonting, i hvarje drag i
sitt uttrycksfulla ansigte. Vidare de kolade bjelkarne, de larmande
soldaterna och bönderna, och öfver hela denna tafla månen med dess
bleka, dallrande sken -- allt detta bildade, säga vi, en högst
egendomlig tafla, tyvärr alls icke främmande för kriget.

"Pojke, du är alldeles galen", ropade Ollola och ämnade just springa
fram, för att, om så behöfdes, med våld rycka sonen från Pekkas sida.
Men han hade knappt tagit ut ett par steg, förrän han såg Rietu,
träffad i bakre delen af hufvudet af en kolfstöt, störta till marken.
Ollola ilade fram och kastade sig på knä vid sonens till utseendet
liflösa kropp.

"Var lugn, gamle Ollola", sade en af bönderna, "slaget var inte så
farligt; pojken kommer sig nog. Den der dufningen gjorde honom godt."

I och med Rietus fall förlorade Pekka helt och hållet det smula mod han
kunnat tilltvinga sig. Men såsom det ofta händer med dylika naturer som
Pekkas, de slå lätt öfver från den ena ytterligheten till den andra. Så
här också. När Pekka nu såg, att han stod ensam och öfvergifven af
alla, brann raseriet i hans själ, och han försökte med all makt att
slita sina bojor, men detta var förgäfves.

"Gå bort, gå bort!" skrek han, när ett par soldater kommo med en snara,
och ögonen voro nära att tränga ut ur sina hålor. "Jag _vill_ inte dö
nu! Tag allt hvad jag eger, men låt mig lefva. Jag ber er derom... Ha,
ni skratta åt min bön. Sätt er bara sjelfva i min ställning, så få ni
väl känna huru det smakar... Nej, tag bort snaran! Hu-u! Tag bort den!"

"Nej, du usle förrädare", dundrade ett par stämmor, "du skall bums in i
evigheten. Gör din bön nu! Fem minuter har du på dig."

Men hurudan var väl den bön, som gick öfver Pirrtiainens skälfvande
läppar? Icke var den sådan, som den borde vara. Han _kunde_ icke bedja
rätt, ty raseriet och den hopplösa förtviflan hade helt och hållet
bemäktigat sig honom.

Innan han visste ordet af, var han kullslagen. En förfärlig ed bröt
fram öfver hans läppar; snaran drogs till och i ett af de högsta träden
på Pirrtiainens gård hängde nu den fordom så högmodige Pekka. Blott ett
par konvulsiviska ryckningar, och allt var slut.

"Vi komma för sent", utbrast Adlercreutz, som med sitt följe nu kom
till ruinerna på samma gång som Elli från sidan störtade fram. "Det var
det jag fruktade, att bönderna skulle tillämpa lynchlagen."

Ett anskri bröt fram öfver den arma Ellis läppar, när hon upptäckte
faderns kropp. Hennes förfäran ökades ännu mera, då hon varseblef
Rietu. Det var nu slut med hennes krafter. Sakta sjönk hon ned öfver
den älskades kropp och förlorade sansen.

"Det var ett allt för hårdt straff", sade Adlercreutz till bönderna.

"Nej, det var alls inte för hårdt", svarade Ollola frimodigt. "Han var
en förrädare, och de äro inte värda någon annan lön."

Generalen teg, ty sanningen i gamle Ollolas ord var obestridlig.

Snart randades en ny tid för Finland. Det blef ryckt ifrån oss, men
friden hägnar nu dessa bygder. Pirrtis uppbyggdes af Rietu, som med sin
hustru Elli der framlefde ett lyckligt lif. Men aldrig glömde Rietu att
för sina barn omtala det sorgliga öde, som drabbat Pekka Pirrtiainen.

"Barn", sade han och pekade på det stora trädet, i hvilket Pekka
blifvit hängd, och som länge stod qvar, "när I sen detta väldiga träd,
så bed Gud bevara er från att blifva fosterlandsförrädare, _ty en sådan
är värd icke blott sina medmenniskors förakt, utan äfven det svåraste
timliga straff man kan upptänka_."